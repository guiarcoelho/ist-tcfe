* NGSPICE simulation script
* BJT amp with feedback
*
* forces current values to be saved
.options savecurrents

.INCLUDE data_sim4.txt
.INCLUDE dataic.txt
*.ic v(6)=8.573530 v(8)=0
.end
.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-6 20e-3

hardcopy transv5vs.ps v(6) v(1)
echo transv5vs_FIG

quit
