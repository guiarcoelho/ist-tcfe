* NGSPICE simulation script
*
* forces current values to be saved
.options savecurrents


.INCLUDE data_sim5.txt
.INCLUDE dataic.txt
*.ic v(6)=8.573530 v(8)=0
* falta automatizar esta merda aqui de cima 
.end
.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

echo "********************************************"
echo  "Frequency analysis"
echo "********************************************"

ac dec 1000 0.1 1MEG

hardcopy acm.ps db(v(6)) db(v(6)-v(8)) db(v(1))
echo acm_FIG

Let phase_v(6) = 180/PI * ph(v(6))
Let phase_v(1) = 180/PI * ph(v(1))
Let phase_v(c) = 180/PI * ph(v(6)-v(8))

hardcopy phase.ps phase_v(6) phase_v(1) phase_v(c)
echo phase_FIG

quit
.endc
